library ieee;
use ieee.std_logic_1164.all;
use work.NbitRegDecs.all;
use work.newBalanceDecs.all;
use work.spinwheelDecs.all;
use work.winDetectorDecs.all;
use work.binToBCDDecs.all;
use work.BCDto7segDecs.all;

use ieee.numeric_std.all; 

entity roulette_top is
  port(SW : in std_logic_vector(17 downto 0);
       KEY : in std_logic_vector(3 downto 0);
       CLOCK_27 : in std_logic;
  		   HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7 : out std_logic_vector(6 downto 0);
  		   LEDG : out std_logic_vector(7 downto 0));
end roulette_top;

architecture impl of roulette_top is
  --wires
  signal spin_result : std_logic_vector(5 downto 0) := "000000";
  signal spin_result_latched : std_logic_vector(5 downto 0) := "000000";
  
  signal money : std_logic_vector(11 downto 0) := "000000000000";
  signal new_money : unsigned(11 downto 0) := "000000000000";
  signal toMoneyFF : unsigned(11 downto 0) := "000000000000";
  
  signal bet1_value : std_logic_vector(5 downto 0) := "000000";
  signal bet2_colour : std_logic_vector(0 downto 0) := "0";
  signal bet2_colour_bit : std_logic := '0';
  signal bet3_dozen : std_logic_vector(1 downto 0) := "00";
    
  signal bet1_wins, bet2_wins, bet3_wins : std_logic := '0';
  
  signal bet1_amt, bet2_amt, bet3_amt : std_logic_vector(2 downto 0) := "000";
  signal bet1_amount, bet2_amount, bet3_amount : unsigned(2 downto 0) := "000";
  
  signal currMoneyBCD : std_logic_vector(11 downto 0);
  signal currMoneyHex : std_logic_vector(20 downto 0); 
  
  signal spinResultBCD : std_logic_vector(7 downto 0);
  signal spinResultHex : std_logic_vector(13 downto 0);

begin
  
  --logic blocks
  num_draw : spinwheel port map(clk => CLOCK_27, rst => KEY(0), spin_result => spin_result);
  
  balance : newBalance port map(money => unsigned(money), new_money => new_money,
            bet1_wins => bet1_wins, bet2_wins => bet2_wins, bet3_wins => bet3_wins,
            bet1_amt => bet1_amount, bet2_amt => bet2_amount, bet3_amt => bet3_amount);
  
  winDetector : win port map(spin_result => unsigned(spin_result),
                 bet1_value => unsigned(bet1_value), bet2_colour => bet2_colour_bit, bet3_dozen => unsigned(bet3_dozen),
                 bet1_wins => bet1_wins, bet2_wins => bet2_wins, bet3_wins => bet3_wins);
  
  --flip flops and conversions
  StateFFspin : NbitReg generic map (6) --spinwheel number
                  port map(rst => KEY(1), clk => KEY(3), D => spin_result, Q => spin_result_latched);
  
  StateFFbetnum : NbitReg generic map (6) --bet number
                  port map(rst => KEY(1), clk => KEY(3), D => SW(8 downto 3), Q => bet1_value);
 
  StateFFbetcolour : NbitReg generic map (1) --bet colour
                  port map(rst => KEY(1), clk => KEY(3), D => SW(12 downto 12), Q => bet2_colour);
  bet2_colour_bit <= bet2_colour(0);
  
  StateFFbetdozen : NbitReg generic map (2) --bet dozen
                  port map(rst => KEY(1), clk => KEY(3), D => SW(17 downto 16), Q => bet3_dozen);
  
  StateFFbet1amt : NbitReg generic map (3) --bet 1 amount
                  port map(rst => KEY(1), clk => KEY(3), D => SW(2 downto 0), Q => bet1_amt);
  
  bet1_amount <= unsigned(bet1_amt);
  
  StateFFbet2amt : NbitReg generic map (3) --bet 2 amount
                  port map(rst => KEY(1), clk => KEY(3), D => SW(11 downto 9), Q => bet2_amt);
  
  bet2_amount <= unsigned(bet2_amt);

  StateFFbet3amt : NbitReg generic map (3) --bet 3 amount
                  port map(rst => KEY(1), clk => KEY(3), D => SW(15 downto 13), Q => bet3_amt);
  
  bet3_amount <= unsigned(bet3_amt);
  
  StateFFmoney : NbitReg generic map (6) --previous money
                  port map(rst => KEY(1), clk => KEY(3), D => std_logic_vector(new_money), Q => money);
  
  toMoneyFF <= unsigned(money);
  
  currMoneyBinToBCD : binToBCD generic map(outDigits => 3, inBits => new_money'LENGTH)
                                  port map(bin => std_logic_vector(new_money), bcd => currMoneyBCD);
                                    
  
  currMoneyBCDTo7Seg :  BCDto7seg generic map(n => 3)
                                        port map(bcd => currMoneyBCD, hex => currMoneyHex); 
  
  spinResultBinToBCD : binToBCD generic map(outDigits => 2, inBits => 6)
                                    port map(bin => std_logic_vector(spin_result), bcd => currMoneyBCD);

  spinResultsBCDToHex : BCDto7seg generic map(n => 2)
                                    port map(bcd => currMoneyBCD, hex => spinResultHex);
                                      
                                                                     
  HEX0 <= currMoneyHex(6 downto 0);
  HEX1 <= currMoneyHex(13 downto 7);
  HEX2 <= currMoneyHex(20 downto 14);

  HEX6 <= spinResultHex(6 downto 0);
  HEX7 <= spinResultHex(13 downto 7);
  
  
  
  LEDG(0) <= bet1_wins;
  LEDG(1) <= bet2_wins;
  LEDG(2) <= bet3_wins;
  
  
  
  
  
  
  
end impl;